// Verilog test fixture created from schematic C:\Users\JaSzw\OneDrive\Pulpit\ISE\Laby4poda\Laby4poda.sch - Sun Apr 05 21:36:02 2020

`timescale 1ns / 1ps

module Laby4poda_Laby4poda_sch_tb();

// Inputs

// Output

// Bidirs

// Instantiate the UUT
   Laby4poda UUT (
		
   );
// Initialize Inputs
   `ifdef auto_init
       initial begin
   `endif
endmodule

`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    10:30:41 04/22/2020 
// Design Name: 
// Module Name:    Laby7sumator_tb 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module Laby7sumator_tb(
input[1:0] a,
input [1:0] b,
output[2:0] y
    );
assign y=a+b;

endmodule

// Verilog test fixture created from schematic C:\Users\JaSzw\OneDrive\Pulpit\ISE\zad2_laby2\zad2.sch - Wed Mar 25 11:29:57 2020

`timescale 1ns / 1ps

module zad2_zad2_sch_tb();

// Inputs

// Output

// Bidirs

// Instantiate the UUT
   zad2 UUT (
		
   );
// Initialize Inputs
   `ifdef auto_init
       initial begin
   `endif
endmodule
